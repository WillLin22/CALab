// this file is to write testbench for module/submodule to check its correctness
`include "cache.vh"
`include "csr_defines.vh"
module WrAligntest ();
    
endmodule