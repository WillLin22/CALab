`define TAGR 20:1
`define VR   0

`define TAGVLEN 21 
`define TAGLEN 20
`define INDEXLEN 8
`define OFFSETLEN 4

`define WAY 2
`define INDEX 256
`define WIDTH 16

`define VATAGR 31:12
`define VAIDXR 11:4
`define VAOFFR 3:0